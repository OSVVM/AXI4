--
--  File Name:         TbAxi4_AlertLogIDManager.vhd
--  Design Unit Name:  Architecture of TestCtrl
--  Revision:          OSVVM MODELS STANDARD VERSION
--
--  Maintainer:        Jim Lewis      email:  jim@synthworks.com
--  Contributor(s):
--     Jim Lewis      jim@synthworks.com
--
--
--  Description:
--      Test transaction source
--
--
--  Developed by:
--        SynthWorks Design Inc.
--        VHDL Training Classes
--        http://www.SynthWorks.com
--
--  Revision History:
--    Date      Version    Description
--    12/2020   2020.12    Initial revision
--
--
--  This file is part of OSVVM.
--  
--  Copyright (c) 2017 - 2021 by SynthWorks Design Inc.  
--  
--  Licensed under the Apache License, Version 2.0 (the "License");
--  you may not use this file except in compliance with the License.
--  You may obtain a copy of the License at
--  
--      https://www.apache.org/licenses/LICENSE-2.0
--  
--  Unless required by applicable law or agreed to in writing, software
--  distributed under the License is distributed on an "AS IS" BASIS,
--  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
--  See the License for the specific language governing permissions and
--  limitations under the License.
--  

architecture AlertLogIDManager of TestCtrl is

  signal TestDone, Sync : integer_barrier := 1 ;
  signal TbManagerID, TbSubordinateID : AlertLogIDType ; 
 
begin

  ------------------------------------------------------------
  -- ControlProc
  --   Set up AlertLog and wait for end of test
  ------------------------------------------------------------
  ControlProc : process
  begin
    -- Initialization of test
    SetTestName("TbAxi4_AlertLogIDManager") ;
    TbManagerID     <= GetAlertLogID("Manager") ;
    TbSubordinateID  <= GetAlertLogID("Subordinate") ;
    SetLogEnable(PASSED, TRUE) ;    -- Enable PASSED logs
    SetLogEnable(INFO, TRUE) ;    -- Enable INFO logs
    SetAlertStopCount(FAILURE, 2) ;    -- Enable INFO logs

    -- Wait for testbench initialization 
    wait for 0 ns ;  wait for 0 ns ;
    TranscriptOpen ;
    SetTranscriptMirror(TRUE) ; 

    -- Wait for Design Reset
    wait until nReset = '1' ;  
    ClearAlerts ;

    -- Wait for test to finish
    WaitForBarrier(TestDone, 35 ms) ;
    AlertIf(now >= 35 ms, "Test finished due to timeout") ;
--    AlertIf(GetAffirmCount < 1, "Test is not Self-Checking");
    
    
    TranscriptClose ; 
    -- Printing differs in different simulators due to differences in process order execution
    -- AffirmIfTranscriptsMatch(PATH_TO_VALIDATED_RESULTS) ;

    EndOfTestReports(ExternalErrors => (FAILURE => -1, ERROR => -1, WARNING => -1)) ; 
    std.env.stop ;
    wait ; 
  end process ControlProc ; 

  ------------------------------------------------------------
  -- ManagerProc
  --   Generate transactions for AxiManager
  ------------------------------------------------------------
  ManagerProc : process
    variable AlertLogID : AlertLogIDType ; 
    variable Count1, Count2 : integer ; 
  begin
    wait until nReset = '1' ;  
    WaitForClock(ManagerRec, 2) ; 
    
    GetAlertLogID(ManagerRec, AlertLogID) ;
    GetErrorCount(ManagerRec, Count1) ;
    AffirmIfEqual(TbManagerID, Count1, 0, "GetErrorCount") ;
    Count2 := GetAlertCount(AlertLogID) ;
    AffirmIfEqual(TbManagerID, Count2, 0, "GetAlertCount") ;
    
    Alert(AlertLogID, "Injected Error 1", ERROR) ;
    GetErrorCount(ManagerRec, Count1) ;
    AffirmIfEqual(TbManagerID, Count1, 1, "GetErrorCount") ;
    Count2 := GetAlertCount(AlertLogID) ;
    AffirmIfEqual(TbManagerID, Count2, 1, "GetAlertCount") ;

    SetAlertStopCount(AlertLogID, FAILURE, 10) ;
    Alert(AlertLogID, "Injected FAILURE 1", FAILURE) ;
    GetErrorCount(ManagerRec, Count1) ;
    AffirmIfEqual(TbManagerID, Count1, 2, "GetErrorCount") ;
    Count2 := GetAlertCount(AlertLogID) ;
    AffirmIfEqual(TbManagerID, Count2, 2, "GetAlertCount") ;

    Alert(AlertLogID, "Injected WARNING 1", WARNING) ;
    GetErrorCount(ManagerRec, Count1) ;
    AffirmIfEqual(TbManagerID, Count1, 3, "GetErrorCount") ;
    Count2 := GetAlertCount(AlertLogID) ;
    AffirmIfEqual(TbManagerID, Count2, 3, "GetAlertCount") ;
    
    WaitForBarrier(TestDone) ;
    wait ;
  end process ManagerProc ;


  ------------------------------------------------------------
  -- SubordinateProc
  --   Generate transactions for AxiSubordinate
  ------------------------------------------------------------
  SubordinateProc : process
    variable Addr : std_logic_vector(AXI_ADDR_WIDTH-1 downto 0) ;
    variable Data : std_logic_vector(AXI_DATA_WIDTH-1 downto 0) ;    
  begin
    wait until nReset = '1' ;  
    WaitForClock(SubordinateRec, 2) ; 
    
    WaitForBarrier(TestDone) ;
    wait ;
  end process SubordinateProc ;


end AlertLogIDManager ;

Configuration TbAxi4_AlertLogIDManager of TbAxi4 is
  for TestHarness
    for TestCtrl_1 : TestCtrl
      use entity work.TestCtrl(AlertLogIDManager) ; 
    end for ; 
  end for ; 
end TbAxi4_AlertLogIDManager ; 