--
--  File Name:         TbAxi4Lite_BasicReadWrite.vhd
--  Design Unit Name:  Architecture of TestCtrl
--  Revision:          OSVVM MODELS STANDARD VERSION
--
--  Maintainer:        Jim Lewis      email:  jim@synthworks.com
--  Contributor(s):
--     Jim Lewis      jim@synthworks.com
--
--
--  Description:
--      Test transaction source
--
--
--  Developed by:
--        SynthWorks Design Inc.
--        VHDL Training Classes
--        http://www.SynthWorks.com
--
--  Revision History:
--    Date       Version    Description
--    09/2017:   2017       Initial revision
--
--
-- Copyright 2017 SynthWorks Design Inc
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
--
architecture BasicReadWrite of TestCtrl is

  signal TestDone : integer_barrier := 1 ;
  constant AXI_ADDR_WIDTH : integer := 32 ; 
  constant AXI_DATA_WIDTH : integer := 32 ; 
 
begin

  ------------------------------------------------------------
  -- ControlProc
  --   Set up AlertLog and wait for end of test
  ------------------------------------------------------------
  ControlProc : process
  begin
    -- Initialization of test
    SetAlertLogName("TbAxi4Lite_BasicReadWrite") ;
    SetLogEnable(PASSED, TRUE) ;    -- Enable PASSED logs
    SetLogEnable(INFO, TRUE) ;    -- Enable INFO logs

    -- Wait for testbench initialization 
    wait for 0 ns ;  wait for 0 ns ;
--    TranscriptOpen("./results/TbAxi4Lite_BasicReadWrite.txt") ;
--    SetTranscriptMirror(TRUE) ; 

    -- Wait for Design Reset
    wait until nReset = '1' ;  
    ClearAlerts ;

    -- Wait for test to finish
    WaitForBarrier(TestDone, 35 ms) ;
    AlertIf(now >= 35 ms, "Test finished due to timeout") ;
    AlertIf(GetAffirmCount < 1, "Test is not Self-Checking");
    
    
--    TranscriptClose ; 
--    AlertIfDiff("./results/TbAxi4Lite_BasicReadWrite.txt", "../sim_shared/validated_results/TbAxi4Lite_BasicReadWrite.txt", "") ; 
    
    print("") ;
    ReportAlerts ; 
    print("") ;
    std.env.stop ; 
    wait ; 
  end process ControlProc ; 

  ------------------------------------------------------------
  -- AxiMasterProc
  --   Generate transactions for AxiMaster
  ------------------------------------------------------------
  AxiMasterProc : process
    variable Data : std_logic_vector(AXI_DATA_WIDTH-1 downto 0) ;
  begin
    wait until nReset = '1' ;  
    NoOp(AxiMasterTransRec, 2) ; 
    log("Write and Read with ByteAddr = 0, 4 Bytes") ;
    MasterWrite(AxiMasterTransRec, X"AAAA_AAA0", X"5555_5555" ) ;
    MasterRead(AxiMasterTransRec,  X"1111_1110", Data) ;
    AffirmIfEqual(Data, X"2222_2222", "Master Read Data: ") ;
    
    log("Write and Read with 1 Byte, and ByteAddr = 0, 1, 2, 3") ; 
    MasterWrite(AxiMasterTransRec, X"AAAA_AAA0", X"11" ) ;
    MasterWrite(AxiMasterTransRec, X"AAAA_AAA1", X"22" ) ;
    MasterWrite(AxiMasterTransRec, X"AAAA_AAA2", X"33" ) ;
    MasterWrite(AxiMasterTransRec, X"AAAA_AAA3", X"44" ) ;
    
    MasterRead(AxiMasterTransRec,  X"1111_1110", Data(7 downto 0)) ;
    AffirmIfEqual(Data(7 downto 0), X"AA", "Master Read Data: ") ;
    MasterRead(AxiMasterTransRec,  X"1111_1111", Data(7 downto 0)) ;
    AffirmIfEqual(Data(7 downto 0), X"BB", "Master Read Data: ") ;
    MasterRead(AxiMasterTransRec,  X"1111_1112", Data(7 downto 0)) ;
    AffirmIfEqual(Data(7 downto 0), X"CC", "Master Read Data: ") ;
    MasterRead(AxiMasterTransRec,  X"1111_1113", Data(7 downto 0)) ;
    AffirmIfEqual(Data(7 downto 0), X"DD", "Master Read Data: ") ;

    log("Write and Read with 2 Bytes, and ByteAddr = 0, 1, 2") ;
    MasterWrite(AxiMasterTransRec, X"BBBB_BBB0", X"2211" ) ;
    MasterWrite(AxiMasterTransRec, X"BBBB_BBB1", X"33_22" ) ;
    MasterWrite(AxiMasterTransRec, X"BBBB_BBB2", X"4433" ) ;

    MasterRead(AxiMasterTransRec,  X"1111_1110", Data(15 downto 0)) ;
    AffirmIfEqual(Data(15 downto 0), X"BBAA", "Master Read Data: ") ;
    MasterRead(AxiMasterTransRec,  X"1111_1111", Data(15 downto 0)) ;
    AffirmIfEqual(Data(15 downto 0), X"CCBB", "Master Read Data: ") ;
    MasterRead(AxiMasterTransRec,  X"1111_1112", Data(15 downto 0)) ;
    AffirmIfEqual(Data(15 downto 0), X"DDCC", "Master Read Data: ") ;

    log("Write and Read with 3 Bytes and ByteAddr = 0. 1") ;
    MasterWrite(AxiMasterTransRec, X"CCCC_CCC0", X"33_2211" ) ;
    MasterWrite(AxiMasterTransRec, X"CCCC_CCC1", X"4433_22" ) ;

    MasterRead(AxiMasterTransRec,  X"1111_1110", Data(23 downto 0)) ;
    AffirmIfEqual(Data(23 downto 0), X"CC_BBAA", "Master Read Data: ") ;
    MasterRead(AxiMasterTransRec,  X"1111_1111", Data(23 downto 0)) ;
    AffirmIfEqual(Data(23 downto 0), X"DDCC_BB", "Master Read Data: ") ;
    
    -- Wait for outputs to propagate and signal TestDone
    NoOp(AxiMasterTransRec, 2) ;
    WaitForBarrier(TestDone) ;
    wait ;
  end process AxiMasterProc ;


  ------------------------------------------------------------
  -- AxiSlaveProc
  --   Generate transactions for AxiSlave
  ------------------------------------------------------------
  AxiSlaveProc : process
    variable Addr : std_logic_vector(AXI_ADDR_WIDTH-1 downto 0) ;
    variable Data : std_logic_vector(AXI_DATA_WIDTH-1 downto 0) ;    
  begin
    NoOp(AxiSlaveTransRec, 2) ; 
    -- Write and Read with ByteAddr = 0, 4 Bytes
    SlaveGetWrite(AxiSlaveTransRec, Addr, Data) ;
    AffirmIfEqual(Addr, X"AAAA_AAA0", "Slave Write Addr: ") ;
    AffirmIfEqual(Data, X"5555_5555", "Slave Write Data: ") ;
    
    SlaveRead(AxiSlaveTransRec, Addr, X"2222_2222") ; 
    AffirmIfEqual(Addr, X"1111_1110", "Slave Read Addr: ") ;

    
    -- Write and Read with 1 Byte, and ByteAddr = 0, 1, 2, 3
    -- MasterWrite(AxiMasterTransRec, X"AAAA_AAA0", X"11" ) ;
    SlaveGetWrite(AxiSlaveTransRec, Addr, Data) ;
    AffirmIfEqual(Addr, X"AAAA_AAA0", "Slave Write Addr: ") ;
    AffirmIfEqual(Data, X"0000_0011", "Slave Write Data: ") ;
    -- MasterWrite(AxiMasterTransRec, X"AAAA_AAA1", X"22" ) ;
    SlaveGetWrite(AxiSlaveTransRec, Addr, Data) ;
    AffirmIfEqual(Addr, X"AAAA_AAA1", "Slave Write Addr: ") ;
    AffirmIfEqual(Data, X"0000_2200", "Slave Write Data: ") ;
    -- MasterWrite(AxiMasterTransRec, X"AAAA_AAA2", X"33" ) ;
    SlaveGetWrite(AxiSlaveTransRec, Addr, Data) ;
    AffirmIfEqual(Addr, X"AAAA_AAA2", "Slave Write Addr: ") ;
    AffirmIfEqual(Data, X"0033_0000", "Slave Write Data: ") ;
    -- MasterWrite(AxiMasterTransRec, X"AAAA_AAA3", X"44" ) ;
    SlaveGetWrite(AxiSlaveTransRec, Addr, Data) ;
    AffirmIfEqual(Addr, X"AAAA_AAA3", "Slave Write Addr: ") ;
    AffirmIfEqual(Data, X"4400_0000", "Slave Write Data: ") ;

    SlaveRead(AxiSlaveTransRec, Addr, X"0000_00AA") ; 
    AffirmIfEqual(Addr, X"1111_1110", "Slave Read Addr: ") ;
    SlaveRead(AxiSlaveTransRec, Addr, X"0000_BB00") ; 
    AffirmIfEqual(Addr, X"1111_1111", "Slave Read Addr: ") ;
    SlaveRead(AxiSlaveTransRec, Addr, X"00CC_0000") ; 
    AffirmIfEqual(Addr, X"1111_1112", "Slave Read Addr: ") ;
    SlaveRead(AxiSlaveTransRec, Addr, X"DD00_0000") ; 
    AffirmIfEqual(Addr, X"1111_1113", "Slave Read Addr: ") ;


    -- Write and Read with 2 Bytes, and ByteAddr = 0, 1, 2
    -- MasterWrite(AxiMasterTransRec, X"BBBB_BBB0", X"2211" ) ;
    SlaveGetWrite(AxiSlaveTransRec, Addr, Data) ;
    AffirmIfEqual(Addr, X"BBBB_BBB0", "Slave Write Addr: ") ;
    AffirmIfEqual(Data, X"0000_2211", "Slave Write Data: ") ;
    -- MasterWrite(AxiMasterTransRec, X"BBBB_BBB1", X"3322" ) ;
    SlaveGetWrite(AxiSlaveTransRec, Addr, Data) ;
    AffirmIfEqual(Addr, X"BBBB_BBB1", "Slave Write Addr: ") ;
    AffirmIfEqual(Data, X"0033_2200", "Slave Write Data: ") ;
    -- MasterWrite(AxiMasterTransRec, X"BBBB_BBB2", X"4433" ) ;
    SlaveGetWrite(AxiSlaveTransRec, Addr, Data) ;
    AffirmIfEqual(Addr, X"BBBB_BBB2", "Slave Write Addr: ") ;
    AffirmIfEqual(Data, X"4433_0000", "Slave Write Data: ") ;

    SlaveRead(AxiSlaveTransRec, Addr, X"0000_BBAA") ; 
    AffirmIfEqual(Addr, X"1111_1110", "Slave Read Addr: ") ;
    SlaveRead(AxiSlaveTransRec, Addr, X"00CC_BB00") ; 
    AffirmIfEqual(Addr, X"1111_1111", "Slave Read Addr: ") ;
    SlaveRead(AxiSlaveTransRec, Addr, X"DDCC_0000") ; 
    AffirmIfEqual(Addr, X"1111_1112", "Slave Read Addr: ") ;

    -- Write and Read with 3 Bytes and ByteAddr = 0. 1
    -- MasterWrite(AxiMasterTransRec, X"CCCC_CCC0", X"332211" ) ;
    SlaveGetWrite(AxiSlaveTransRec, Addr, Data) ;
    AffirmIfEqual(Addr, X"CCCC_CCC0", "Slave Write Addr: ") ;
    AffirmIfEqual(Data, X"0033_2211", "Slave Write Data: ") ;
    -- MasterWrite(AxiMasterTransRec, X"CCCC_CCC1", X"443322" ) ;
    SlaveGetWrite(AxiSlaveTransRec, Addr, Data) ;
    AffirmIfEqual(Addr, X"CCCC_CCC1", "Slave Write Addr: ") ;
    AffirmIfEqual(Data, X"4433_2200", "Slave Write Data: ") ;

    SlaveRead(AxiSlaveTransRec, Addr, X"00CC_BBAA") ; 
    AffirmIfEqual(Addr, X"1111_1110", "Slave Read Addr: ") ;
    SlaveRead(AxiSlaveTransRec, Addr, X"DDCC_BB00") ; 
    AffirmIfEqual(Addr, X"1111_1111", "Slave Read Addr: ") ;


    -- Wait for outputs to propagate and signal TestDone
    NoOp(AxiSlaveTransRec, 2) ;
    WaitForBarrier(TestDone) ;
    wait ;
  end process AxiSlaveProc ;


end BasicReadWrite ;

Configuration TbAxi4Lite_BasicReadWrite of TbAxi4Lite is
  for TestHarness
    for TestCtrl_1 : TestCtrl
      use entity work.TestCtrl(BasicReadWrite) ; 
    end for ; 
  end for ; 
end TbAxi4Lite_BasicReadWrite ; 